module ConvolutionUnit (
    parameter DATA_WIDTH = 32;
    parameter KERNEL_SIZE = 3;
    parameter

    input clk, reset;
    input []
);
    
endmodule